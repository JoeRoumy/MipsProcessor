module test();

main Main();

endmodule

